@80000000
6F 00 80 04 73 2F 20 34 93 0F 80 00 63 08 FF 03
93 0F 90 00 63 04 FF 03 93 0F B0 00 63 00 FF 03
13 0F 00 00 63 04 0F 00 67 00 0F 00 73 2F 20 34
63 54 0F 00 6F 00 40 00 93 E1 91 53 17 1F 00 00
23 22 3F FC 6F F0 9F FF 93 00 00 00 13 01 00 00
93 01 00 00 13 02 00 00 93 02 00 00 13 03 00 00
93 03 00 00 13 04 00 00 93 04 00 00 13 05 00 00
93 05 00 00 13 06 00 00 93 06 00 00 13 07 00 00
93 07 00 00 13 08 00 00 93 08 00 00 13 09 00 00
93 09 00 00 13 0A 00 00 93 0A 00 00 13 0B 00 00
93 0B 00 00 13 0C 00 00 93 0C 00 00 13 0D 00 00
93 0D 00 00 13 0E 00 00 93 0E 00 00 13 0F 00 00
93 0F 00 00 73 25 40 F1 63 10 05 00 97 02 00 00
93 82 02 01 73 90 52 30 73 50 00 18 97 02 00 00
93 82 02 02 73 90 52 30 B7 02 00 80 93 82 F2 FF
73 90 02 3B 93 02 F0 01 73 90 02 3A 73 50 40 30
97 02 00 00 93 82 42 01 73 90 52 30 73 50 20 30
73 50 30 30 93 01 00 00 97 02 00 00 93 82 C2 EE
73 90 52 30 13 05 10 00 13 15 F5 01 63 4C 05 00
0F 00 F0 0F 93 01 10 00 93 08 D0 05 13 05 00 00
73 00 00 00 93 02 00 00 63 8A 02 00 73 90 52 10
B7 B2 00 00 93 82 92 10 73 90 22 30 73 50 00 30
97 02 00 00 93 82 42 01 73 90 12 34 73 25 40 F1
73 00 20 30 93 01 20 00 93 00 00 00 13 01 00 00
63 D6 20 00 63 18 30 30 63 16 30 00 E3 DE 20 FE
63 12 30 30 93 01 30 00 93 00 10 00 13 01 10 00
63 D6 20 00 63 18 30 2E 63 16 30 00 E3 DE 20 FE
63 12 30 2E 93 01 40 00 93 00 F0 FF 13 01 F0 FF
63 D6 20 00 63 18 30 2C 63 16 30 00 E3 DE 20 FE
63 12 30 2C 93 01 50 00 93 00 10 00 13 01 00 00
63 D6 20 00 63 18 30 2A 63 16 30 00 E3 DE 20 FE
63 12 30 2A 93 01 60 00 93 00 10 00 13 01 F0 FF
63 D6 20 00 63 18 30 28 63 16 30 00 E3 DE 20 FE
63 12 30 28 93 01 70 00 93 00 F0 FF 13 01 E0 FF
63 D6 20 00 63 18 30 26 63 16 30 00 E3 DE 20 FE
63 12 30 26 93 01 80 00 93 00 00 00 13 01 10 00
63 D4 20 00 63 14 30 00 63 16 30 24 E3 DE 20 FE
93 01 90 00 93 00 F0 FF 13 01 10 00 63 D4 20 00
63 14 30 00 63 18 30 22 E3 DE 20 FE 93 01 A0 00
93 00 E0 FF 13 01 F0 FF 63 D4 20 00 63 14 30 00
63 1A 30 20 E3 DE 20 FE 93 01 B0 00 93 00 E0 FF
13 01 10 00 63 D4 20 00 63 14 30 00 63 1C 30 1E
E3 DE 20 FE 93 01 C0 00 13 02 00 00 93 00 F0 FF
13 01 00 00 63 D0 20 1E 13 02 12 00 93 02 20 00
E3 16 52 FE 93 01 D0 00 13 02 00 00 93 00 F0 FF
13 01 00 00 13 00 00 00 63 DE 20 1A 13 02 12 00
93 02 20 00 E3 14 52 FE 93 01 E0 00 13 02 00 00
93 00 F0 FF 13 01 00 00 13 00 00 00 13 00 00 00
63 DA 20 18 13 02 12 00 93 02 20 00 E3 12 52 FE
93 01 F0 00 13 02 00 00 93 00 F0 FF 13 00 00 00
13 01 00 00 63 D8 20 16 13 02 12 00 93 02 20 00
E3 14 52 FE 93 01 00 01 13 02 00 00 93 00 F0 FF
13 00 00 00 13 01 00 00 13 00 00 00 63 D4 20 14
13 02 12 00 93 02 20 00 E3 12 52 FE 93 01 10 01
13 02 00 00 93 00 F0 FF 13 00 00 00 13 00 00 00
13 01 00 00 63 D0 20 12 13 02 12 00 93 02 20 00
E3 12 52 FE 93 01 20 01 13 02 00 00 93 00 F0 FF
13 01 00 00 63 D0 20 10 13 02 12 00 93 02 20 00
E3 16 52 FE 93 01 30 01 13 02 00 00 93 00 F0 FF
13 01 00 00 13 00 00 00 63 DE 20 0C 13 02 12 00
93 02 20 00 E3 14 52 FE 93 01 40 01 13 02 00 00
93 00 F0 FF 13 01 00 00 13 00 00 00 13 00 00 00
63 DA 20 0A 13 02 12 00 93 02 20 00 E3 12 52 FE
93 01 50 01 13 02 00 00 93 00 F0 FF 13 00 00 00
13 01 00 00 63 D8 20 08 13 02 12 00 93 02 20 00
E3 14 52 FE 93 01 60 01 13 02 00 00 93 00 F0 FF
13 00 00 00 13 01 00 00 13 00 00 00 63 D4 20 06
13 02 12 00 93 02 20 00 E3 12 52 FE 93 01 70 01
13 02 00 00 93 00 F0 FF 13 00 00 00 13 00 00 00
13 01 00 00 63 D0 20 04 13 02 12 00 93 02 20 00
E3 12 52 FE 93 00 10 00 63 DA 00 00 93 80 10 00
93 80 10 00 93 80 10 00 93 80 10 00 93 80 10 00
93 80 10 00 93 03 30 00 93 01 80 01 63 94 70 00
63 10 30 02 0F 00 F0 0F 63 80 01 00 93 91 11 00
93 E1 11 00 93 08 D0 05 13 85 01 00 73 00 00 00
0F 00 F0 0F 93 01 10 00 93 08 D0 05 13 05 00 00
73 00 00 00 73 10 00 C0 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00
@80001000
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00
