@80000000
6F 00 80 04 73 2F 20 34 93 0F 80 00 63 08 FF 03
93 0F 90 00 63 04 FF 03 93 0F B0 00 63 00 FF 03
13 0F 00 00 63 04 0F 00 67 00 0F 00 73 2F 20 34
63 54 0F 00 6F 00 40 00 93 E1 91 53 17 1F 00 00
23 22 3F FC 6F F0 9F FF 93 00 00 00 13 01 00 00
93 01 00 00 13 02 00 00 93 02 00 00 13 03 00 00
93 03 00 00 13 04 00 00 93 04 00 00 13 05 00 00
93 05 00 00 13 06 00 00 93 06 00 00 13 07 00 00
93 07 00 00 13 08 00 00 93 08 00 00 13 09 00 00
93 09 00 00 13 0A 00 00 93 0A 00 00 13 0B 00 00
93 0B 00 00 13 0C 00 00 93 0C 00 00 13 0D 00 00
93 0D 00 00 13 0E 00 00 93 0E 00 00 13 0F 00 00
93 0F 00 00 73 25 40 F1 63 10 05 00 97 02 00 00
93 82 02 01 73 90 52 30 73 50 00 18 97 02 00 00
93 82 02 02 73 90 52 30 B7 02 00 80 93 82 F2 FF
73 90 02 3B 93 02 F0 01 73 90 02 3A 73 50 40 30
97 02 00 00 93 82 42 01 73 90 52 30 73 50 20 30
73 50 30 30 93 01 00 00 97 02 00 00 93 82 C2 EE
73 90 52 30 13 05 10 00 13 15 F5 01 63 4C 05 00
0F 00 F0 0F 93 01 10 00 93 08 D0 05 13 05 00 00
73 00 00 00 93 02 00 00 63 8A 02 00 73 90 52 10
B7 B2 00 00 93 82 92 10 73 90 22 30 73 50 00 30
97 02 00 00 93 82 42 01 73 90 12 34 73 25 40 F1
73 00 20 30 93 01 20 00 93 02 00 00 17 03 00 00
13 03 03 01 E7 02 03 00 6F 00 00 0E 17 03 00 00
13 03 C3 FF 63 9A 62 0C 93 01 30 00 97 02 00 00
93 82 02 01 E7 82 02 00 6F 00 00 0C 17 03 00 00
13 03 C3 FF 63 9A 62 0A 93 01 40 00 13 02 00 00
17 03 00 00 13 03 03 01 E7 06 03 00 63 1E 30 08
13 02 12 00 93 02 20 00 E3 14 52 FE 93 01 50 00
13 02 00 00 17 03 00 00 13 03 43 01 13 00 00 00
E7 06 03 00 63 1A 30 06 13 02 12 00 93 02 20 00
E3 12 52 FE 93 01 60 00 13 02 00 00 17 03 00 00
13 03 83 01 13 00 00 00 13 00 00 00 E7 06 03 00
63 14 30 04 13 02 12 00 93 02 20 00 E3 10 52 FE
93 02 10 00 17 03 00 00 13 03 C3 01 67 00 C3 FF
93 82 12 00 93 82 12 00 93 82 12 00 93 82 12 00
93 82 12 00 93 82 12 00 93 03 40 00 93 01 70 00
63 94 72 00 63 10 30 02 0F 00 F0 0F 63 80 01 00
93 91 11 00 93 E1 11 00 93 08 D0 05 13 85 01 00
73 00 00 00 0F 00 F0 0F 93 01 10 00 93 08 D0 05
13 05 00 00 73 00 00 00 73 10 00 C0 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00
@80001000
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00
