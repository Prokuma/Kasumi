@80000000
6F 00 80 04 73 2F 20 34 93 0F 80 00 63 08 FF 03
93 0F 90 00 63 04 FF 03 93 0F B0 00 63 00 FF 03
13 0F 00 00 63 04 0F 00 67 00 0F 00 73 2F 20 34
63 54 0F 00 6F 00 40 00 93 E1 91 53 17 1F 00 00
23 22 3F FC 6F F0 9F FF 93 00 00 00 13 01 00 00
93 01 00 00 13 02 00 00 93 02 00 00 13 03 00 00
93 03 00 00 13 04 00 00 93 04 00 00 13 05 00 00
93 05 00 00 13 06 00 00 93 06 00 00 13 07 00 00
93 07 00 00 13 08 00 00 93 08 00 00 13 09 00 00
93 09 00 00 13 0A 00 00 93 0A 00 00 13 0B 00 00
93 0B 00 00 13 0C 00 00 93 0C 00 00 13 0D 00 00
93 0D 00 00 13 0E 00 00 93 0E 00 00 13 0F 00 00
93 0F 00 00 73 25 40 F1 63 10 05 00 97 02 00 00
93 82 02 01 73 90 52 30 73 50 00 18 97 02 00 00
93 82 02 02 73 90 52 30 B7 02 00 80 93 82 F2 FF
73 90 02 3B 93 02 F0 01 73 90 02 3A 73 50 40 30
97 02 00 00 93 82 42 01 73 90 52 30 73 50 20 30
73 50 30 30 93 01 00 00 97 02 00 00 93 82 C2 EE
73 90 52 30 13 05 10 00 13 15 F5 01 63 4C 05 00
0F 00 F0 0F 93 01 10 00 93 08 D0 05 13 05 00 00
73 00 00 00 93 02 00 00 63 8A 02 00 73 90 52 10
B7 B2 00 00 93 82 92 10 73 90 22 30 73 50 00 30
97 02 00 00 93 82 42 01 73 90 12 34 73 25 40 F1
73 00 20 30 97 20 00 00 93 80 C0 E8 13 01 A0 0A
23 90 20 00 03 97 00 00 93 03 A0 0A 93 01 20 00
63 1E 77 44 97 20 00 00 93 80 C0 E6 37 B1 FF FF
13 01 01 A0 23 91 20 00 03 97 20 00 B7 B3 FF FF
93 83 03 A0 93 01 30 00 63 1A 77 42 97 20 00 00
93 80 40 E4 37 11 EF BE 13 01 01 AA 23 92 20 00
03 A7 40 00 B7 13 EF BE 93 83 03 AA 93 01 40 00
63 16 77 40 97 20 00 00 93 80 C0 E1 37 A1 FF FF
13 01 A1 00 23 93 20 00 03 97 60 00 B7 A3 FF FF
93 83 A3 00 93 01 50 00 63 12 77 3E 97 20 00 00
93 80 20 E0 13 01 A0 0A 23 9D 20 FE 03 97 A0 FF
93 03 A0 0A 93 01 60 00 63 12 77 3C 97 20 00 00
93 80 20 DE 37 B1 FF FF 13 01 01 A0 23 9E 20 FE
03 97 C0 FF B7 B3 FF FF 93 83 03 A0 93 01 70 00
63 1E 77 38 97 20 00 00 93 80 A0 DB 37 11 00 00
13 01 01 AA 23 9F 20 FE 03 97 E0 FF B7 13 00 00
93 83 03 AA 93 01 80 00 63 1A 77 36 97 20 00 00
93 80 20 D9 37 A1 FF FF 13 01 A1 00 23 90 20 00
03 97 00 00 B7 A3 FF FF 93 83 A3 00 93 01 90 00
63 16 77 34 97 20 00 00 93 80 C0 D6 37 51 34 12
13 01 81 67 13 82 00 FE 23 10 22 02 83 92 00 00
B7 53 00 00 93 83 83 67 93 01 A0 00 63 90 72 32
97 20 00 00 93 80 00 D4 37 31 00 00 13 01 81 09
93 80 B0 FF A3 93 20 00 17 22 00 00 13 02 A2 D2
83 12 02 00 B7 33 00 00 93 83 83 09 93 01 B0 00
63 96 72 2E 93 01 C0 00 13 02 00 00 B7 D0 FF FF
93 80 D0 CD 17 21 00 00 13 01 C1 CE 23 10 11 00
03 17 01 00 B7 D3 FF FF 93 83 D3 CD 63 10 77 2C
13 02 12 00 93 02 20 00 E3 1A 52 FC 93 01 D0 00
13 02 00 00 B7 C0 FF FF 93 80 D0 CC 17 21 00 00
13 01 41 CB 13 00 00 00 23 11 11 00 03 17 21 00
B7 C3 FF FF 93 83 D3 CC 63 12 77 28 13 02 12 00
93 02 20 00 E3 18 52 FC 93 01 E0 00 13 02 00 00
B7 C0 FF FF 93 80 C0 BC 17 21 00 00 13 01 81 C7
13 00 00 00 13 00 00 00 23 12 11 00 03 17 41 00
B7 C3 FF FF 93 83 C3 BC 63 12 77 24 13 02 12 00
93 02 20 00 E3 16 52 FC 93 01 F0 00 13 02 00 00
B7 B0 FF FF 93 80 C0 BB 13 00 00 00 17 21 00 00
13 01 41 C3 23 13 11 00 03 17 61 00 B7 B3 FF FF
93 83 C3 BB 63 14 77 20 13 02 12 00 93 02 20 00
E3 18 52 FC 93 01 00 01 13 02 00 00 B7 B0 FF FF
93 80 B0 AB 13 00 00 00 17 21 00 00 13 01 81 BF
13 00 00 00 23 14 11 00 03 17 81 00 B7 B3 FF FF
93 83 B3 AB 63 14 77 1C 13 02 12 00 93 02 20 00
E3 16 52 FC 93 01 10 01 13 02 00 00 B7 E0 FF FF
93 80 B0 AA 13 00 00 00 13 00 00 00 17 21 00 00
13 01 41 BB 23 15 11 00 03 17 A1 00 B7 E3 FF FF
93 83 B3 AA 63 14 77 18 13 02 12 00 93 02 20 00
E3 16 52 FC 93 01 20 01 13 02 00 00 17 21 00 00
13 01 41 B8 B7 20 00 00 93 80 30 23 23 10 11 00
03 17 01 00 B7 23 00 00 93 83 33 23 63 18 77 14
13 02 12 00 93 02 20 00 E3 1A 52 FC 93 01 30 01
13 02 00 00 17 21 00 00 13 01 C1 B4 B7 10 00 00
93 80 30 22 13 00 00 00 23 11 11 00 03 17 21 00
B7 13 00 00 93 83 33 22 63 1A 77 10 13 02 12 00
93 02 20 00 E3 18 52 FC 93 01 40 01 13 02 00 00
17 21 00 00 13 01 01 B1 B7 10 00 00 93 80 20 12
13 00 00 00 13 00 00 00 23 12 11 00 03 17 41 00
B7 13 00 00 93 83 23 12 63 1A 77 0C 13 02 12 00
93 02 20 00 E3 16 52 FC 93 01 50 01 13 02 00 00
17 21 00 00 13 01 01 AD 13 00 00 00 93 00 20 11
23 13 11 00 03 17 61 00 93 03 20 11 63 10 77 0A
13 02 12 00 93 02 20 00 E3 1C 52 FC 93 01 60 01
13 02 00 00 17 21 00 00 13 01 C1 A9 13 00 00 00
93 00 10 01 13 00 00 00 23 14 11 00 03 17 81 00
93 03 10 01 63 14 77 06 13 02 12 00 93 02 20 00
E3 1A 52 FC 93 01 70 01 13 02 00 00 17 21 00 00
13 01 41 A6 13 00 00 00 13 00 00 00 B7 30 00 00
93 80 10 00 23 15 11 00 03 17 A1 00 B7 33 00 00
93 83 13 00 63 14 77 02 13 02 12 00 93 02 20 00
E3 16 52 FC 37 C5 00 00 13 05 F5 EE 97 25 00 00
93 85 45 A2 23 93 A5 00 63 10 30 02 0F 00 F0 0F
63 80 01 00 93 91 11 00 93 E1 11 00 93 08 D0 05
13 85 01 00 73 00 00 00 0F 00 F0 0F 93 01 10 00
93 08 D0 05 13 05 00 00 73 00 00 00 73 10 00 C0
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00
@80001000
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00
@80002000
EF BE EF BE EF BE EF BE EF BE EF BE EF BE EF BE
EF BE EF BE 00 00 00 00 00 00 00 00 00 00 00 00
