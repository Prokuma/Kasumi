@80000000
6F 00 80 04 73 2F 20 34 93 0F 80 00 63 08 FF 03
93 0F 90 00 63 04 FF 03 93 0F B0 00 63 00 FF 03
13 0F 00 00 63 04 0F 00 67 00 0F 00 73 2F 20 34
63 54 0F 00 6F 00 40 00 93 E1 91 53 17 1F 00 00
23 22 3F FC 6F F0 9F FF 93 00 00 00 13 01 00 00
93 01 00 00 13 02 00 00 93 02 00 00 13 03 00 00
93 03 00 00 13 04 00 00 93 04 00 00 13 05 00 00
93 05 00 00 13 06 00 00 93 06 00 00 13 07 00 00
93 07 00 00 13 08 00 00 93 08 00 00 13 09 00 00
93 09 00 00 13 0A 00 00 93 0A 00 00 13 0B 00 00
93 0B 00 00 13 0C 00 00 93 0C 00 00 13 0D 00 00
93 0D 00 00 13 0E 00 00 93 0E 00 00 13 0F 00 00
93 0F 00 00 73 25 40 F1 63 10 05 00 97 02 00 00
93 82 02 01 73 90 52 30 73 50 00 18 97 02 00 00
93 82 02 02 73 90 52 30 B7 02 00 80 93 82 F2 FF
73 90 02 3B 93 02 F0 01 73 90 02 3A 73 50 40 30
97 02 00 00 93 82 42 01 73 90 52 30 73 50 20 30
73 50 30 30 93 01 00 00 97 02 00 00 93 82 C2 EE
73 90 52 30 13 05 10 00 13 15 F5 01 63 4C 05 00
0F 00 F0 0F 93 01 10 00 93 08 D0 05 13 05 00 00
73 00 00 00 93 02 00 00 63 8A 02 00 73 90 52 10
B7 B2 00 00 93 82 92 10 73 90 22 30 73 50 00 30
97 02 00 00 93 82 42 01 73 90 12 34 73 25 40 F1
73 00 20 30 97 20 00 00 93 80 C0 E8 03 A7 00 00
B7 03 FF 00 93 83 F3 0F 93 01 20 00 63 1A 77 26
97 20 00 00 93 80 00 E7 03 A7 40 00 B7 03 01 FF
93 83 03 F0 93 01 30 00 63 1C 77 24 97 20 00 00
93 80 40 E5 03 A7 80 00 B7 13 F0 0F 93 83 03 FF
93 01 40 00 63 1E 77 22 97 20 00 00 93 80 80 E3
03 A7 C0 00 B7 F3 0F F0 93 83 F3 00 93 01 50 00
63 10 77 22 97 20 00 00 93 80 80 E2 03 A7 40 FF
B7 03 FF 00 93 83 F3 0F 93 01 60 00 63 12 77 20
97 20 00 00 93 80 C0 E0 03 A7 80 FF B7 03 01 FF
93 83 03 F0 93 01 70 00 63 14 77 1E 97 20 00 00
93 80 00 DF 03 A7 C0 FF B7 13 F0 0F 93 83 03 FF
93 01 80 00 63 16 77 1C 97 20 00 00 93 80 40 DD
03 A7 00 00 B7 F3 0F F0 93 83 F3 00 93 01 90 00
63 18 77 1A 97 20 00 00 93 80 C0 DA 93 80 00 FE
83 A2 00 02 B7 03 FF 00 93 83 F3 0F 93 01 A0 00
63 98 72 18 97 20 00 00 93 80 C0 D8 93 80 D0 FF
83 A2 70 00 B7 03 01 FF 93 83 03 F0 93 01 B0 00
63 98 72 16 93 01 C0 00 13 02 00 00 97 20 00 00
93 80 80 D6 03 A7 40 00 13 03 07 00 B7 13 F0 0F
93 83 03 FF 63 16 73 14 13 02 12 00 93 02 20 00
E3 1E 52 FC 93 01 D0 00 13 02 00 00 97 20 00 00
93 80 C0 D3 03 A7 40 00 13 00 00 00 13 03 07 00
B7 F3 0F F0 93 83 F3 00 63 1C 73 10 13 02 12 00
93 02 20 00 E3 1C 52 FC 93 01 E0 00 13 02 00 00
97 20 00 00 93 80 00 D0 03 A7 40 00 13 00 00 00
13 00 00 00 13 03 07 00 B7 03 01 FF 93 83 03 F0
63 10 73 0E 13 02 12 00 93 02 20 00 E3 1A 52 FC
93 01 F0 00 13 02 00 00 97 20 00 00 93 80 C0 CC
03 A7 40 00 B7 13 F0 0F 93 83 03 FF 63 1A 77 0A
13 02 12 00 93 02 20 00 E3 10 52 FE 93 01 00 01
13 02 00 00 97 20 00 00 93 80 40 CA 13 00 00 00
03 A7 40 00 B7 F3 0F F0 93 83 F3 00 63 12 77 08
13 02 12 00 93 02 20 00 E3 1E 52 FC 93 01 10 01
13 02 00 00 97 20 00 00 93 80 C0 C6 13 00 00 00
13 00 00 00 03 A7 40 00 B7 03 01 FF 93 83 03 F0
63 18 77 04 13 02 12 00 93 02 20 00 E3 1C 52 FC
97 22 00 00 93 82 02 C4 03 A1 02 00 13 01 20 00
93 03 20 00 93 01 20 01 63 14 71 02 97 22 00 00
93 82 42 C2 03 A1 02 00 13 00 00 00 13 01 20 00
93 03 20 00 93 01 30 01 63 14 71 00 63 10 30 02
0F 00 F0 0F 63 80 01 00 93 91 11 00 93 E1 11 00
93 08 D0 05 13 85 01 00 73 00 00 00 0F 00 F0 0F
93 01 10 00 93 08 D0 05 13 05 00 00 73 00 00 00
73 10 00 C0 00 00 00 00 00 00 00 00
@80001000
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00
@80002000
FF 00 FF 00 00 FF 00 FF F0 0F F0 0F 0F F0 0F F0
