@80000000
6F 00 80 04 73 2F 20 34 93 0F 80 00 63 08 FF 03
93 0F 90 00 63 04 FF 03 93 0F B0 00 63 00 FF 03
13 0F 00 00 63 04 0F 00 67 00 0F 00 73 2F 20 34
63 54 0F 00 6F 00 40 00 93 E1 91 53 17 1F 00 00
23 22 3F FC 6F F0 9F FF 93 00 00 00 13 01 00 00
93 01 00 00 13 02 00 00 93 02 00 00 13 03 00 00
93 03 00 00 13 04 00 00 93 04 00 00 13 05 00 00
93 05 00 00 13 06 00 00 93 06 00 00 13 07 00 00
93 07 00 00 13 08 00 00 93 08 00 00 13 09 00 00
93 09 00 00 13 0A 00 00 93 0A 00 00 13 0B 00 00
93 0B 00 00 13 0C 00 00 93 0C 00 00 13 0D 00 00
93 0D 00 00 13 0E 00 00 93 0E 00 00 13 0F 00 00
93 0F 00 00 73 25 40 F1 63 10 05 00 97 02 00 00
93 82 02 01 73 90 52 30 73 50 00 18 97 02 00 00
93 82 02 02 73 90 52 30 B7 02 00 80 93 82 F2 FF
73 90 02 3B 93 02 F0 01 73 90 02 3A 73 50 40 30
97 02 00 00 93 82 42 01 73 90 52 30 73 50 20 30
73 50 30 30 93 01 00 00 97 02 00 00 93 82 C2 EE
73 90 52 30 13 05 10 00 13 15 F5 01 63 4C 05 00
0F 00 F0 0F 93 01 10 00 93 08 D0 05 13 05 00 00
73 00 00 00 93 02 00 00 63 8A 02 00 73 90 52 10
B7 B2 00 00 93 82 92 10 73 90 22 30 73 50 00 30
97 02 00 00 93 82 42 01 73 90 12 34 73 25 40 F1
73 00 20 30 97 20 00 00 93 80 C0 E8 13 01 A0 FA
23 80 20 00 03 87 00 00 93 03 A0 FA 93 01 20 00
63 1C 77 3C 97 20 00 00 93 80 C0 E6 13 01 00 00
A3 80 20 00 03 87 10 00 93 03 00 00 93 01 30 00
63 1C 77 3A 97 20 00 00 93 80 C0 E4 37 F1 FF FF
13 01 01 FA 23 81 20 00 03 97 20 00 B7 F3 FF FF
93 83 03 FA 93 01 40 00 63 18 77 38 97 20 00 00
93 80 40 E2 13 01 A0 00 A3 81 20 00 03 87 30 00
93 03 A0 00 93 01 50 00 63 18 77 36 97 20 00 00
93 80 B0 E0 13 01 A0 FA A3 8E 20 FE 03 87 D0 FF
93 03 A0 FA 93 01 60 00 63 18 77 34 97 20 00 00
93 80 B0 DE 13 01 00 00 23 8F 20 FE 03 87 E0 FF
93 03 00 00 93 01 70 00 63 18 77 32 97 20 00 00
93 80 B0 DC 13 01 00 FA A3 8F 20 FE 03 87 F0 FF
93 03 00 FA 93 01 80 00 63 18 77 30 97 20 00 00
93 80 B0 DA 13 01 A0 00 23 80 20 00 03 87 00 00
93 03 A0 00 93 01 90 00 63 18 77 2E 97 20 00 00
93 80 C0 D8 37 51 34 12 13 01 81 67 13 82 00 FE
23 00 22 02 83 82 00 00 93 03 80 07 93 01 A0 00
63 94 72 2C 97 20 00 00 93 80 40 D6 37 31 00 00
13 01 81 09 93 80 A0 FF A3 83 20 00 17 22 00 00
13 02 D2 D4 83 02 02 00 93 03 80 F9 93 01 B0 00
63 9C 72 28 93 01 C0 00 13 02 00 00 93 00 D0 FD
17 21 00 00 13 01 01 D2 23 00 11 00 03 07 01 00
93 03 D0 FD 63 1A 77 26 13 02 12 00 93 02 20 00
E3 1E 52 FC 93 01 D0 00 13 02 00 00 93 00 D0 FC
17 21 00 00 13 01 01 CF 13 00 00 00 A3 00 11 00
03 07 11 00 93 03 D0 FC 63 10 77 24 13 02 12 00
93 02 20 00 E3 1C 52 FC 93 01 E0 00 13 02 00 00
93 00 C0 FC 17 21 00 00 13 01 C1 CB 13 00 00 00
13 00 00 00 23 01 11 00 03 07 21 00 93 03 C0 FC
63 14 77 20 13 02 12 00 93 02 20 00 E3 1A 52 FC
93 01 F0 00 13 02 00 00 93 00 C0 FB 13 00 00 00
17 21 00 00 13 01 01 C8 A3 01 11 00 03 07 31 00
93 03 C0 FB 63 1A 77 1C 13 02 12 00 93 02 20 00
E3 1C 52 FC 93 01 00 01 13 02 00 00 93 00 B0 FB
13 00 00 00 17 21 00 00 13 01 C1 C4 13 00 00 00
23 02 11 00 03 07 41 00 93 03 B0 FB 63 1E 77 18
13 02 12 00 93 02 20 00 E3 1A 52 FC 93 01 10 01
13 02 00 00 93 00 B0 FA 13 00 00 00 13 00 00 00
17 21 00 00 13 01 01 C1 A3 02 11 00 03 07 51 00
93 03 B0 FA 63 12 77 16 13 02 12 00 93 02 20 00
E3 1A 52 FC 93 01 20 01 13 02 00 00 17 21 00 00
13 01 41 BE 93 00 30 03 23 00 11 00 03 07 01 00
93 03 30 03 63 1A 77 12 13 02 12 00 93 02 20 00
E3 1E 52 FC 93 01 30 01 13 02 00 00 17 21 00 00
13 01 41 BB 93 00 30 02 13 00 00 00 A3 00 11 00
03 07 11 00 93 03 30 02 63 10 77 10 13 02 12 00
93 02 20 00 E3 1C 52 FC 93 01 40 01 13 02 00 00
17 21 00 00 13 01 01 B8 93 00 20 02 13 00 00 00
13 00 00 00 23 01 11 00 03 07 21 00 93 03 20 02
63 14 77 0C 13 02 12 00 93 02 20 00 E3 1A 52 FC
93 01 50 01 13 02 00 00 17 21 00 00 13 01 81 B4
13 00 00 00 93 00 20 01 A3 01 11 00 03 07 31 00
93 03 20 01 63 1A 77 08 13 02 12 00 93 02 20 00
E3 1C 52 FC 93 01 60 01 13 02 00 00 17 21 00 00
13 01 41 B1 13 00 00 00 93 00 10 01 13 00 00 00
23 02 11 00 03 07 41 00 93 03 10 01 63 1E 77 04
13 02 12 00 93 02 20 00 E3 1A 52 FC 93 01 70 01
13 02 00 00 17 21 00 00 13 01 C1 AD 13 00 00 00
13 00 00 00 93 00 10 00 A3 02 11 00 03 07 51 00
93 03 10 00 63 12 77 02 13 02 12 00 93 02 20 00
E3 1A 52 FC 13 05 F0 0E 97 25 00 00 93 85 85 AA
A3 81 A5 00 63 10 30 02 0F 00 F0 0F 63 80 01 00
93 91 11 00 93 E1 11 00 93 08 D0 05 13 85 01 00
73 00 00 00 0F 00 F0 0F 93 01 10 00 93 08 D0 05
13 05 00 00 73 00 00 00 73 10 00 C0 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00
@80001000
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00
@80002000
EF EF EF EF EF EF EF EF EF EF 00 00 00 00 00 00
